`timescale 1ns/1ns
`include "encoder.v"

module encoder_tb;

    reg [3:0] bcd;
    wire [6:0] Y;

    encoder teste(bcd,Y);
    
    initial begin
        $dumpfile("encoder.vcd");
        $dumpvars(0, encoder_tb);

        bcd = 4'b0000; #10;
        bcd = 4'b0001; #10;
        bcd = 4'b0010; #10;
        bcd = 4'b0011; #10;
        bcd = 4'b0100; #10;
        bcd = 4'b0101; #10;
        bcd = 4'b0110; #10;
        bcd = 4'b0111; #10;
        bcd = 4'b1000; #10;
        bcd = 4'b1001; #10;
        bcd = 4'b1010; #10;
        bcd = 4'b1011; #10;
        bcd = 4'b1100; #10;
        bcd = 4'b1101; #10;
        bcd = 4'b1110; #10;
        bcd = 4'b1111; #10;

        $display("Teste completo");
    end

endmodule